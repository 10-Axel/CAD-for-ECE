
.MODEL NMOS NMOS (                                LEVEL   = 7
+ TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 2.3549E17      VTH0    = 0.3750766
+K1      = 0.5842025      K2      = 1.245202E-3    K3      = 1E-3
+K3B     = 0.0295587      W0      = 1E-7           NLX     = 1.597846E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 1.3022984      DVT1    = 0.4021873      DVT2    = 7.631374E-3
+U0      = 296.8451012    UA      = -1.179955E-9   UB      = 2.32616E-18
+UC      = 7.593301E-11   VSAT    = 1.747147E5     A0      = 2
+AGS     = 0.452647       B0      = 5.506962E-8    B1      = 2.640458E-6
+KETA    = -6.860244E-3   A1      = 7.885522E-4    A2      = 0.3119338
+RDSW    = 105            PRWG    = 0.4826         PRWB    = -0.2
+WR      = 1              WINT    = 4.410779E-9    LINT    = 2.045919E-8
+XL      = 0              XW      = -1E-8          DWG     = -2.610453E-9
+DWB     = -4.344942E-9   VOFF    = -0.0948017     NFACTOR = 2.1860065
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 1.991317E-3    ETAB    = 6.028975E-5
+DSUB    = 0.0217897      PCLM    = 1.7062594      PDIBLC1 = 0.2320546
+PDIBLC2 = 1.670588E-3    PDIBLCB = -0.1           DROUT   = 0.8388608
+PSCBE1  = 1.904263E10    PSCBE2  = 1.546939E-8    PVAG    = 0
+DELTA   = 0.01           RSH     = 7.1            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 6.7E-10        CGSO    = 6.7E-10        CGBO    = 1E-12
+CJ      = 9.550345E-4    PB      = 0.8            MJ      = 0.3762949
+CJSW    = 2.083251E-10   PBSW    = 0.8            MJSW    = 0.1269477
+CJSWG   = 3.3E-10        PBSWG   = 0.8            MJSWG   = 0.1269477
+CF      = 0              PVTH0   = -2.369258E-3   PRDSW   = -1.2091688
+PK2     = 1.845281E-3    WKETA   = -2.040084E-3   LKETA   = -1.266704E-3
+PU0     = 1.0932981      PUA     = -2.56934E-11   PUB     = 0
+PVSAT   = 2E3            PETA0   = 1E-4           PKETA   = -3.350276E-3    )
*
.MODEL PMOS PMOS (                                LEVEL   = 7
+ TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 4.1589E17      VTH0    = -0.3936726
+K1      = 0.5750728      K2      = 0.0235926      K3      = 0.1590089
+K3B     = 4.2687016      W0      = 1E-6           NLX     = 1.033999E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.5560978      DVT1    = 0.2490116      DVT2    = 0.1
+U0      = 112.5106786    UA      = 1.45072E-9     UB      = 1.195045E-21
+UC      = -1E-10         VSAT    = 1.168535E5     A0      = 1.7211984
+AGS     = 0.3806925      B0      = 4.296252E-7    B1      = 1.288698E-6
+KETA    = 0.0201833      A1      = 0.2328472      A2      = 0.3
+RDSW    = 198.7483291    PRWG    = 0.5            PRWB    = -0.4971827
+WR      = 1              WINT    = 0              LINT    = 2.943206E-8
+XL      = 0              XW      = -1E-8          DWG     = -1.949253E-8
+DWB     = -2.824041E-9   VOFF    = -0.0979832     NFACTOR = 1.9624066
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 7.282772E-4    ETAB    = -3.818572E-4
+DSUB    = 1.518344E-3    PCLM    = 1.4728931      PDIBLC1 = 2.138043E-3
+PDIBLC2 = -9.966066E-6   PDIBLCB = -1E-3          DROUT   = 4.276128E-4
+PSCBE1  = 4.850167E10    PSCBE2  = 5E-10          PVAG    = 0
+DELTA   = 0.01           RSH     = 8.2            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 7.47E-10       CGSO    = 7.47E-10       CGBO    = 1E-12
+CJ      = 1.180017E-3    PB      = 0.8560642      MJ      = 0.4146818
+CJSW    = 2.046463E-10   PBSW    = 0.9123142      MJSW    = 0.316175
+CJSWG   = 4.22E-10       PBSWG   = 0.9123142      MJSWG   = 0.316175
+CF      = 0              PVTH0   = 8.456598E-4    PRDSW   = 8.4838247
+PK2     = 1.338191E-3    WKETA   = 0.0246885      LKETA   = -2.016897E-3
+PU0     = -1.5089586     PUA     = -5.51646E-11   PUB     = 1E-21
+PVSAT   = 50             PETA0   = 1E-4           PKETA   = -3.316832E-3    )

.subckt INVERTER Ni No
Mn No Ni 0 0 NMOS W=0.18u L=0.19u
Mp No Ni Ndd Ndd PMOS W=0.45u L=0.18u
Vdd Ndd 0 dc 1.8v
.ends
X1 N1 No1 INVERTER
X2 No1 No2 INVERTER
M1 Ndi Nclk N1 N1 NMOS  W=0.9u L=0.18u
M2 No2 Nclkb N1 N1 NMOS W=0.9u L=0.18u
Vi Ndi 0 pulse(0 1.8v 1u 0 1n 10u  20u)
Vclk Nclk 0 pulse(0 1.8v 3u 1n 1n 10u 20u)
Vclkb Nclkb 0 pulse(1.8v 0 3u 1n 1n 10u 20u)
.tran 1n 80u
.probe
.end










